// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Feb 18 2018 15:14:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "chip" view "INTERFACE"

module chip (
    PMOD,
    ADR,
    DAT,
    clk,
    RAMWE,
    RAMOE,
    RAMCS);

    output [55:0] PMOD;
    output [18:0] ADR;
    output [15:0] DAT;
    input clk;
    output RAMWE;
    output RAMOE;
    output RAMCS;

    wire N__2714;
    wire N__2713;
    wire N__2712;
    wire N__2703;
    wire N__2702;
    wire N__2701;
    wire N__2694;
    wire N__2693;
    wire N__2692;
    wire N__2685;
    wire N__2684;
    wire N__2683;
    wire N__2676;
    wire N__2675;
    wire N__2674;
    wire N__2667;
    wire N__2666;
    wire N__2665;
    wire N__2658;
    wire N__2657;
    wire N__2656;
    wire N__2649;
    wire N__2648;
    wire N__2647;
    wire N__2640;
    wire N__2639;
    wire N__2638;
    wire N__2631;
    wire N__2630;
    wire N__2629;
    wire N__2622;
    wire N__2621;
    wire N__2620;
    wire N__2613;
    wire N__2612;
    wire N__2611;
    wire N__2604;
    wire N__2603;
    wire N__2602;
    wire N__2595;
    wire N__2594;
    wire N__2593;
    wire N__2586;
    wire N__2585;
    wire N__2584;
    wire N__2577;
    wire N__2576;
    wire N__2575;
    wire N__2568;
    wire N__2567;
    wire N__2566;
    wire N__2559;
    wire N__2558;
    wire N__2557;
    wire N__2550;
    wire N__2549;
    wire N__2548;
    wire N__2541;
    wire N__2540;
    wire N__2539;
    wire N__2532;
    wire N__2531;
    wire N__2530;
    wire N__2523;
    wire N__2522;
    wire N__2521;
    wire N__2514;
    wire N__2513;
    wire N__2512;
    wire N__2505;
    wire N__2504;
    wire N__2503;
    wire N__2496;
    wire N__2495;
    wire N__2494;
    wire N__2487;
    wire N__2486;
    wire N__2485;
    wire N__2478;
    wire N__2477;
    wire N__2476;
    wire N__2469;
    wire N__2468;
    wire N__2467;
    wire N__2460;
    wire N__2459;
    wire N__2458;
    wire N__2451;
    wire N__2450;
    wire N__2449;
    wire N__2442;
    wire N__2441;
    wire N__2440;
    wire N__2433;
    wire N__2432;
    wire N__2431;
    wire N__2424;
    wire N__2423;
    wire N__2422;
    wire N__2415;
    wire N__2414;
    wire N__2413;
    wire N__2406;
    wire N__2405;
    wire N__2404;
    wire N__2397;
    wire N__2396;
    wire N__2395;
    wire N__2388;
    wire N__2387;
    wire N__2386;
    wire N__2379;
    wire N__2378;
    wire N__2377;
    wire N__2370;
    wire N__2369;
    wire N__2368;
    wire N__2361;
    wire N__2360;
    wire N__2359;
    wire N__2352;
    wire N__2351;
    wire N__2350;
    wire N__2343;
    wire N__2342;
    wire N__2341;
    wire N__2334;
    wire N__2333;
    wire N__2332;
    wire N__2325;
    wire N__2324;
    wire N__2323;
    wire N__2316;
    wire N__2315;
    wire N__2314;
    wire N__2307;
    wire N__2306;
    wire N__2305;
    wire N__2298;
    wire N__2297;
    wire N__2296;
    wire N__2289;
    wire N__2288;
    wire N__2287;
    wire N__2280;
    wire N__2279;
    wire N__2278;
    wire N__2271;
    wire N__2270;
    wire N__2269;
    wire N__2262;
    wire N__2261;
    wire N__2260;
    wire N__2253;
    wire N__2252;
    wire N__2251;
    wire N__2244;
    wire N__2243;
    wire N__2242;
    wire N__2235;
    wire N__2234;
    wire N__2233;
    wire N__2226;
    wire N__2225;
    wire N__2224;
    wire N__2217;
    wire N__2216;
    wire N__2215;
    wire N__2208;
    wire N__2207;
    wire N__2206;
    wire N__2199;
    wire N__2198;
    wire N__2197;
    wire N__2190;
    wire N__2189;
    wire N__2188;
    wire N__2181;
    wire N__2180;
    wire N__2179;
    wire N__2172;
    wire N__2171;
    wire N__2170;
    wire N__2163;
    wire N__2162;
    wire N__2161;
    wire N__2154;
    wire N__2153;
    wire N__2152;
    wire N__2145;
    wire N__2144;
    wire N__2143;
    wire N__2136;
    wire N__2135;
    wire N__2134;
    wire N__2127;
    wire N__2126;
    wire N__2125;
    wire N__2118;
    wire N__2117;
    wire N__2116;
    wire N__2109;
    wire N__2108;
    wire N__2107;
    wire N__2100;
    wire N__2099;
    wire N__2098;
    wire N__2091;
    wire N__2090;
    wire N__2089;
    wire N__2082;
    wire N__2081;
    wire N__2080;
    wire N__2073;
    wire N__2072;
    wire N__2071;
    wire N__2064;
    wire N__2063;
    wire N__2062;
    wire N__2055;
    wire N__2054;
    wire N__2053;
    wire N__2046;
    wire N__2045;
    wire N__2044;
    wire N__2037;
    wire N__2036;
    wire N__2035;
    wire N__2028;
    wire N__2027;
    wire N__2026;
    wire N__2019;
    wire N__2018;
    wire N__2017;
    wire N__2010;
    wire N__2009;
    wire N__2008;
    wire N__2001;
    wire N__2000;
    wire N__1999;
    wire N__1992;
    wire N__1991;
    wire N__1990;
    wire N__1983;
    wire N__1982;
    wire N__1981;
    wire N__1974;
    wire N__1973;
    wire N__1972;
    wire N__1965;
    wire N__1964;
    wire N__1963;
    wire N__1956;
    wire N__1955;
    wire N__1954;
    wire N__1947;
    wire N__1946;
    wire N__1945;
    wire N__1938;
    wire N__1937;
    wire N__1936;
    wire N__1929;
    wire N__1928;
    wire N__1927;
    wire N__1920;
    wire N__1919;
    wire N__1918;
    wire N__1911;
    wire N__1910;
    wire N__1909;
    wire N__1902;
    wire N__1901;
    wire N__1900;
    wire N__1893;
    wire N__1892;
    wire N__1891;
    wire N__1884;
    wire N__1883;
    wire N__1882;
    wire N__1875;
    wire N__1874;
    wire N__1873;
    wire N__1866;
    wire N__1865;
    wire N__1864;
    wire N__1847;
    wire N__1846;
    wire N__1843;
    wire N__1840;
    wire N__1835;
    wire N__1832;
    wire N__1831;
    wire N__1828;
    wire N__1825;
    wire N__1820;
    wire N__1817;
    wire N__1816;
    wire N__1813;
    wire N__1810;
    wire N__1805;
    wire N__1802;
    wire N__1801;
    wire N__1798;
    wire N__1795;
    wire N__1792;
    wire N__1789;
    wire N__1784;
    wire N__1781;
    wire N__1778;
    wire N__1775;
    wire N__1772;
    wire N__1769;
    wire N__1766;
    wire N__1763;
    wire N__1760;
    wire N__1757;
    wire N__1754;
    wire N__1751;
    wire N__1748;
    wire N__1745;
    wire N__1742;
    wire N__1739;
    wire N__1736;
    wire N__1733;
    wire N__1730;
    wire N__1727;
    wire N__1724;
    wire N__1721;
    wire N__1718;
    wire N__1715;
    wire N__1712;
    wire N__1709;
    wire N__1706;
    wire N__1703;
    wire N__1700;
    wire N__1697;
    wire N__1694;
    wire N__1691;
    wire N__1690;
    wire N__1689;
    wire N__1688;
    wire N__1679;
    wire N__1676;
    wire N__1673;
    wire N__1670;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1658;
    wire N__1655;
    wire N__1652;
    wire N__1649;
    wire N__1646;
    wire N__1643;
    wire N__1640;
    wire N__1637;
    wire N__1634;
    wire N__1631;
    wire N__1628;
    wire N__1625;
    wire N__1622;
    wire N__1619;
    wire N__1616;
    wire N__1613;
    wire N__1610;
    wire N__1607;
    wire N__1604;
    wire N__1601;
    wire N__1598;
    wire N__1595;
    wire N__1592;
    wire N__1589;
    wire N__1586;
    wire N__1583;
    wire N__1580;
    wire N__1577;
    wire N__1574;
    wire N__1571;
    wire N__1568;
    wire N__1565;
    wire N__1562;
    wire N__1559;
    wire N__1556;
    wire N__1553;
    wire N__1550;
    wire N__1547;
    wire N__1544;
    wire N__1541;
    wire N__1538;
    wire N__1535;
    wire N__1532;
    wire N__1529;
    wire N__1526;
    wire N__1523;
    wire N__1520;
    wire N__1517;
    wire N__1514;
    wire N__1511;
    wire N__1508;
    wire N__1505;
    wire N__1502;
    wire N__1499;
    wire N__1496;
    wire N__1493;
    wire N__1490;
    wire N__1487;
    wire N__1484;
    wire N__1481;
    wire N__1478;
    wire N__1475;
    wire N__1472;
    wire N__1469;
    wire N__1468;
    wire N__1465;
    wire N__1462;
    wire N__1459;
    wire N__1458;
    wire N__1455;
    wire N__1452;
    wire N__1449;
    wire N__1446;
    wire N__1443;
    wire N__1440;
    wire N__1437;
    wire N__1434;
    wire N__1431;
    wire N__1428;
    wire N__1425;
    wire N__1422;
    wire N__1419;
    wire VCCG0;
    wire GNDG0;
    wire CONSTANT_ONE_NET;
    wire \my_alternate.countZ0Z_0 ;
    wire bfn_19_6_0_;
    wire \my_alternate.countZ0Z_1 ;
    wire \my_alternate.count_cry_0 ;
    wire \my_alternate.countZ0Z_2 ;
    wire \my_alternate.count_cry_1 ;
    wire \my_alternate.countZ0Z_3 ;
    wire \my_alternate.count_cry_2 ;
    wire \my_alternate.countZ0Z_4 ;
    wire \my_alternate.count_cry_3 ;
    wire \my_alternate.countZ0Z_5 ;
    wire \my_alternate.count_cry_4 ;
    wire \my_alternate.countZ0Z_6 ;
    wire \my_alternate.count_cry_5 ;
    wire \my_alternate.countZ0Z_7 ;
    wire \my_alternate.count_cry_6 ;
    wire \my_alternate.count_cry_7 ;
    wire \my_alternate.countZ0Z_8 ;
    wire bfn_19_7_0_;
    wire \my_alternate.countZ0Z_9 ;
    wire \my_alternate.count_cry_8 ;
    wire \my_alternate.countZ0Z_10 ;
    wire \my_alternate.count_cry_9 ;
    wire \my_alternate.countZ0Z_11 ;
    wire \my_alternate.count_cry_10 ;
    wire \my_alternate.countZ0Z_12 ;
    wire \my_alternate.count_cry_11 ;
    wire \my_alternate.countZ0Z_13 ;
    wire \my_alternate.count_cry_12 ;
    wire \my_alternate.countZ0Z_14 ;
    wire \my_alternate.count_cry_13 ;
    wire \my_alternate.countZ0Z_15 ;
    wire \my_alternate.count_cry_14 ;
    wire \my_alternate.count_cry_15 ;
    wire \my_alternate.countZ0Z_16 ;
    wire bfn_19_8_0_;
    wire \my_alternate.countZ0Z_17 ;
    wire \my_alternate.count_cry_16 ;
    wire \my_alternate.countZ0Z_18 ;
    wire \my_alternate.count_cry_17 ;
    wire \my_alternate.countZ0Z_19 ;
    wire \my_alternate.count_cry_18 ;
    wire \my_alternate.countZ0Z_20 ;
    wire \my_alternate.count_cry_19 ;
    wire \my_alternate.countZ0Z_21 ;
    wire \my_alternate.count_cry_20 ;
    wire \my_alternate.countZ0Z_22 ;
    wire \my_alternate.count_cry_21 ;
    wire \my_alternate.countZ0Z_23 ;
    wire \my_alternate.count_cry_22 ;
    wire \my_alternate.count_cry_23 ;
    wire bfn_19_9_0_;
    wire clk_c_g;
    wire PMOD_c_52;
    wire PMOD_c_i_52;
    wire _gnd_net_;

    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2712),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__2714),
            .DIN(N__2713),
            .DOUT(N__2712),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__2714),
            .PADOUT(N__2713),
            .PADIN(N__2712),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_0_iopad (
            .OE(N__2703),
            .DIN(N__2702),
            .DOUT(N__2701),
            .PACKAGEPIN(ADR[0]));
    defparam ADR_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_0_preio (
            .PADOEN(N__2703),
            .PADOUT(N__2702),
            .PADIN(N__2701),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_1_iopad (
            .OE(N__2694),
            .DIN(N__2693),
            .DOUT(N__2692),
            .PACKAGEPIN(ADR[1]));
    defparam ADR_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_1_preio (
            .PADOEN(N__2694),
            .PADOUT(N__2693),
            .PADIN(N__2692),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_10_iopad (
            .OE(N__2685),
            .DIN(N__2684),
            .DOUT(N__2683),
            .PACKAGEPIN(ADR[10]));
    defparam ADR_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_10_preio (
            .PADOEN(N__2685),
            .PADOUT(N__2684),
            .PADIN(N__2683),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_11_iopad (
            .OE(N__2676),
            .DIN(N__2675),
            .DOUT(N__2674),
            .PACKAGEPIN(ADR[11]));
    defparam ADR_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_11_preio (
            .PADOEN(N__2676),
            .PADOUT(N__2675),
            .PADIN(N__2674),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_12_iopad (
            .OE(N__2667),
            .DIN(N__2666),
            .DOUT(N__2665),
            .PACKAGEPIN(ADR[12]));
    defparam ADR_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_12_preio (
            .PADOEN(N__2667),
            .PADOUT(N__2666),
            .PADIN(N__2665),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_13_iopad (
            .OE(N__2658),
            .DIN(N__2657),
            .DOUT(N__2656),
            .PACKAGEPIN(ADR[13]));
    defparam ADR_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_13_preio (
            .PADOEN(N__2658),
            .PADOUT(N__2657),
            .PADIN(N__2656),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_14_iopad (
            .OE(N__2649),
            .DIN(N__2648),
            .DOUT(N__2647),
            .PACKAGEPIN(ADR[14]));
    defparam ADR_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_14_preio (
            .PADOEN(N__2649),
            .PADOUT(N__2648),
            .PADIN(N__2647),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_15_iopad (
            .OE(N__2640),
            .DIN(N__2639),
            .DOUT(N__2638),
            .PACKAGEPIN(ADR[15]));
    defparam ADR_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_15_preio (
            .PADOEN(N__2640),
            .PADOUT(N__2639),
            .PADIN(N__2638),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_16_iopad (
            .OE(N__2631),
            .DIN(N__2630),
            .DOUT(N__2629),
            .PACKAGEPIN(ADR[16]));
    defparam ADR_obuf_16_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_16_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_16_preio (
            .PADOEN(N__2631),
            .PADOUT(N__2630),
            .PADIN(N__2629),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_17_iopad (
            .OE(N__2622),
            .DIN(N__2621),
            .DOUT(N__2620),
            .PACKAGEPIN(ADR[17]));
    defparam ADR_obuf_17_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_17_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_17_preio (
            .PADOEN(N__2622),
            .PADOUT(N__2621),
            .PADIN(N__2620),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_18_iopad (
            .OE(N__2613),
            .DIN(N__2612),
            .DOUT(N__2611),
            .PACKAGEPIN(ADR[18]));
    defparam ADR_obuf_18_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_18_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_18_preio (
            .PADOEN(N__2613),
            .PADOUT(N__2612),
            .PADIN(N__2611),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_2_iopad (
            .OE(N__2604),
            .DIN(N__2603),
            .DOUT(N__2602),
            .PACKAGEPIN(ADR[2]));
    defparam ADR_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_2_preio (
            .PADOEN(N__2604),
            .PADOUT(N__2603),
            .PADIN(N__2602),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_3_iopad (
            .OE(N__2595),
            .DIN(N__2594),
            .DOUT(N__2593),
            .PACKAGEPIN(ADR[3]));
    defparam ADR_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_3_preio (
            .PADOEN(N__2595),
            .PADOUT(N__2594),
            .PADIN(N__2593),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_4_iopad (
            .OE(N__2586),
            .DIN(N__2585),
            .DOUT(N__2584),
            .PACKAGEPIN(ADR[4]));
    defparam ADR_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_4_preio (
            .PADOEN(N__2586),
            .PADOUT(N__2585),
            .PADIN(N__2584),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_5_iopad (
            .OE(N__2577),
            .DIN(N__2576),
            .DOUT(N__2575),
            .PACKAGEPIN(ADR[5]));
    defparam ADR_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_5_preio (
            .PADOEN(N__2577),
            .PADOUT(N__2576),
            .PADIN(N__2575),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_6_iopad (
            .OE(N__2568),
            .DIN(N__2567),
            .DOUT(N__2566),
            .PACKAGEPIN(ADR[6]));
    defparam ADR_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_6_preio (
            .PADOEN(N__2568),
            .PADOUT(N__2567),
            .PADIN(N__2566),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_7_iopad (
            .OE(N__2559),
            .DIN(N__2558),
            .DOUT(N__2557),
            .PACKAGEPIN(ADR[7]));
    defparam ADR_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_7_preio (
            .PADOEN(N__2559),
            .PADOUT(N__2558),
            .PADIN(N__2557),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_8_iopad (
            .OE(N__2550),
            .DIN(N__2549),
            .DOUT(N__2548),
            .PACKAGEPIN(ADR[8]));
    defparam ADR_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_8_preio (
            .PADOEN(N__2550),
            .PADOUT(N__2549),
            .PADIN(N__2548),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD ADR_obuf_9_iopad (
            .OE(N__2541),
            .DIN(N__2540),
            .DOUT(N__2539),
            .PACKAGEPIN(ADR[9]));
    defparam ADR_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam ADR_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO ADR_obuf_9_preio (
            .PADOEN(N__2541),
            .PADOUT(N__2540),
            .PADIN(N__2539),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_0_iopad (
            .OE(N__2532),
            .DIN(N__2531),
            .DOUT(N__2530),
            .PACKAGEPIN(DAT[0]));
    defparam DAT_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_0_preio (
            .PADOEN(N__2532),
            .PADOUT(N__2531),
            .PADIN(N__2530),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_1_iopad (
            .OE(N__2523),
            .DIN(N__2522),
            .DOUT(N__2521),
            .PACKAGEPIN(DAT[1]));
    defparam DAT_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_1_preio (
            .PADOEN(N__2523),
            .PADOUT(N__2522),
            .PADIN(N__2521),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_10_iopad (
            .OE(N__2514),
            .DIN(N__2513),
            .DOUT(N__2512),
            .PACKAGEPIN(DAT[10]));
    defparam DAT_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_10_preio (
            .PADOEN(N__2514),
            .PADOUT(N__2513),
            .PADIN(N__2512),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_11_iopad (
            .OE(N__2505),
            .DIN(N__2504),
            .DOUT(N__2503),
            .PACKAGEPIN(DAT[11]));
    defparam DAT_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_11_preio (
            .PADOEN(N__2505),
            .PADOUT(N__2504),
            .PADIN(N__2503),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_12_iopad (
            .OE(N__2496),
            .DIN(N__2495),
            .DOUT(N__2494),
            .PACKAGEPIN(DAT[12]));
    defparam DAT_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_12_preio (
            .PADOEN(N__2496),
            .PADOUT(N__2495),
            .PADIN(N__2494),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_13_iopad (
            .OE(N__2487),
            .DIN(N__2486),
            .DOUT(N__2485),
            .PACKAGEPIN(DAT[13]));
    defparam DAT_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_13_preio (
            .PADOEN(N__2487),
            .PADOUT(N__2486),
            .PADIN(N__2485),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_14_iopad (
            .OE(N__2478),
            .DIN(N__2477),
            .DOUT(N__2476),
            .PACKAGEPIN(DAT[14]));
    defparam DAT_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_14_preio (
            .PADOEN(N__2478),
            .PADOUT(N__2477),
            .PADIN(N__2476),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_15_iopad (
            .OE(N__2469),
            .DIN(N__2468),
            .DOUT(N__2467),
            .PACKAGEPIN(DAT[15]));
    defparam DAT_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_15_preio (
            .PADOEN(N__2469),
            .PADOUT(N__2468),
            .PADIN(N__2467),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_2_iopad (
            .OE(N__2460),
            .DIN(N__2459),
            .DOUT(N__2458),
            .PACKAGEPIN(DAT[2]));
    defparam DAT_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_2_preio (
            .PADOEN(N__2460),
            .PADOUT(N__2459),
            .PADIN(N__2458),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_3_iopad (
            .OE(N__2451),
            .DIN(N__2450),
            .DOUT(N__2449),
            .PACKAGEPIN(DAT[3]));
    defparam DAT_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_3_preio (
            .PADOEN(N__2451),
            .PADOUT(N__2450),
            .PADIN(N__2449),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_4_iopad (
            .OE(N__2442),
            .DIN(N__2441),
            .DOUT(N__2440),
            .PACKAGEPIN(DAT[4]));
    defparam DAT_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_4_preio (
            .PADOEN(N__2442),
            .PADOUT(N__2441),
            .PADIN(N__2440),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_5_iopad (
            .OE(N__2433),
            .DIN(N__2432),
            .DOUT(N__2431),
            .PACKAGEPIN(DAT[5]));
    defparam DAT_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_5_preio (
            .PADOEN(N__2433),
            .PADOUT(N__2432),
            .PADIN(N__2431),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_6_iopad (
            .OE(N__2424),
            .DIN(N__2423),
            .DOUT(N__2422),
            .PACKAGEPIN(DAT[6]));
    defparam DAT_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_6_preio (
            .PADOEN(N__2424),
            .PADOUT(N__2423),
            .PADIN(N__2422),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_7_iopad (
            .OE(N__2415),
            .DIN(N__2414),
            .DOUT(N__2413),
            .PACKAGEPIN(DAT[7]));
    defparam DAT_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_7_preio (
            .PADOEN(N__2415),
            .PADOUT(N__2414),
            .PADIN(N__2413),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_8_iopad (
            .OE(N__2406),
            .DIN(N__2405),
            .DOUT(N__2404),
            .PACKAGEPIN(DAT[8]));
    defparam DAT_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_8_preio (
            .PADOEN(N__2406),
            .PADOUT(N__2405),
            .PADIN(N__2404),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD DAT_obuf_9_iopad (
            .OE(N__2397),
            .DIN(N__2396),
            .DOUT(N__2395),
            .PACKAGEPIN(DAT[9]));
    defparam DAT_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DAT_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO DAT_obuf_9_preio (
            .PADOEN(N__2397),
            .PADOUT(N__2396),
            .PADIN(N__2395),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuf_52_iopad (
            .OE(N__2388),
            .DIN(N__2387),
            .DOUT(N__2386),
            .PACKAGEPIN(PMOD[52]));
    defparam PMOD_obuf_52_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuf_52_preio.PIN_TYPE=6'b011001;
    PRE_IO PMOD_obuf_52_preio (
            .PADOEN(N__2388),
            .PADOUT(N__2387),
            .PADIN(N__2386),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1847),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuf_53_iopad (
            .OE(N__2379),
            .DIN(N__2378),
            .DOUT(N__2377),
            .PACKAGEPIN(PMOD[53]));
    defparam PMOD_obuf_53_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuf_53_preio.PIN_TYPE=6'b011001;
    PRE_IO PMOD_obuf_53_preio (
            .PADOEN(N__2379),
            .PADOUT(N__2378),
            .PADIN(N__2377),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1801),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuf_54_iopad (
            .OE(N__2370),
            .DIN(N__2369),
            .DOUT(N__2368),
            .PACKAGEPIN(PMOD[54]));
    defparam PMOD_obuf_54_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuf_54_preio.PIN_TYPE=6'b011001;
    PRE_IO PMOD_obuf_54_preio (
            .PADOEN(N__2370),
            .PADOUT(N__2369),
            .PADIN(N__2368),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1846),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuf_55_iopad (
            .OE(N__2361),
            .DIN(N__2360),
            .DOUT(N__2359),
            .PACKAGEPIN(PMOD[55]));
    defparam PMOD_obuf_55_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuf_55_preio.PIN_TYPE=6'b011001;
    PRE_IO PMOD_obuf_55_preio (
            .PADOEN(N__2361),
            .PADOUT(N__2360),
            .PADIN(N__2359),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1805),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_0_iopad (
            .OE(N__2352),
            .DIN(N__2351),
            .DOUT(N__2350),
            .PACKAGEPIN(PMOD[0]));
    defparam PMOD_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_0_preio (
            .PADOEN(N__2352),
            .PADOUT(N__2351),
            .PADIN(N__2350),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_1_iopad (
            .OE(N__2343),
            .DIN(N__2342),
            .DOUT(N__2341),
            .PACKAGEPIN(PMOD[1]));
    defparam PMOD_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_1_preio (
            .PADOEN(N__2343),
            .PADOUT(N__2342),
            .PADIN(N__2341),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_10_iopad (
            .OE(N__2334),
            .DIN(N__2333),
            .DOUT(N__2332),
            .PACKAGEPIN(PMOD[10]));
    defparam PMOD_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_10_preio (
            .PADOEN(N__2334),
            .PADOUT(N__2333),
            .PADIN(N__2332),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_11_iopad (
            .OE(N__2325),
            .DIN(N__2324),
            .DOUT(N__2323),
            .PACKAGEPIN(PMOD[11]));
    defparam PMOD_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_11_preio (
            .PADOEN(N__2325),
            .PADOUT(N__2324),
            .PADIN(N__2323),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_12_iopad (
            .OE(N__2316),
            .DIN(N__2315),
            .DOUT(N__2314),
            .PACKAGEPIN(PMOD[12]));
    defparam PMOD_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_12_preio (
            .PADOEN(N__2316),
            .PADOUT(N__2315),
            .PADIN(N__2314),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_13_iopad (
            .OE(N__2307),
            .DIN(N__2306),
            .DOUT(N__2305),
            .PACKAGEPIN(PMOD[13]));
    defparam PMOD_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_13_preio (
            .PADOEN(N__2307),
            .PADOUT(N__2306),
            .PADIN(N__2305),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_14_iopad (
            .OE(N__2298),
            .DIN(N__2297),
            .DOUT(N__2296),
            .PACKAGEPIN(PMOD[14]));
    defparam PMOD_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_14_preio (
            .PADOEN(N__2298),
            .PADOUT(N__2297),
            .PADIN(N__2296),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_15_iopad (
            .OE(N__2289),
            .DIN(N__2288),
            .DOUT(N__2287),
            .PACKAGEPIN(PMOD[15]));
    defparam PMOD_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_15_preio (
            .PADOEN(N__2289),
            .PADOUT(N__2288),
            .PADIN(N__2287),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_16_iopad (
            .OE(N__2280),
            .DIN(N__2279),
            .DOUT(N__2278),
            .PACKAGEPIN(PMOD[16]));
    defparam PMOD_obuft_16_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_16_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_16_preio (
            .PADOEN(N__2280),
            .PADOUT(N__2279),
            .PADIN(N__2278),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_17_iopad (
            .OE(N__2271),
            .DIN(N__2270),
            .DOUT(N__2269),
            .PACKAGEPIN(PMOD[17]));
    defparam PMOD_obuft_17_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_17_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_17_preio (
            .PADOEN(N__2271),
            .PADOUT(N__2270),
            .PADIN(N__2269),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_18_iopad (
            .OE(N__2262),
            .DIN(N__2261),
            .DOUT(N__2260),
            .PACKAGEPIN(PMOD[18]));
    defparam PMOD_obuft_18_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_18_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_18_preio (
            .PADOEN(N__2262),
            .PADOUT(N__2261),
            .PADIN(N__2260),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_19_iopad (
            .OE(N__2253),
            .DIN(N__2252),
            .DOUT(N__2251),
            .PACKAGEPIN(PMOD[19]));
    defparam PMOD_obuft_19_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_19_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_19_preio (
            .PADOEN(N__2253),
            .PADOUT(N__2252),
            .PADIN(N__2251),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_2_iopad (
            .OE(N__2244),
            .DIN(N__2243),
            .DOUT(N__2242),
            .PACKAGEPIN(PMOD[2]));
    defparam PMOD_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_2_preio (
            .PADOEN(N__2244),
            .PADOUT(N__2243),
            .PADIN(N__2242),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_20_iopad (
            .OE(N__2235),
            .DIN(N__2234),
            .DOUT(N__2233),
            .PACKAGEPIN(PMOD[20]));
    defparam PMOD_obuft_20_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_20_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_20_preio (
            .PADOEN(N__2235),
            .PADOUT(N__2234),
            .PADIN(N__2233),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_21_iopad (
            .OE(N__2226),
            .DIN(N__2225),
            .DOUT(N__2224),
            .PACKAGEPIN(PMOD[21]));
    defparam PMOD_obuft_21_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_21_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_21_preio (
            .PADOEN(N__2226),
            .PADOUT(N__2225),
            .PADIN(N__2224),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_22_iopad (
            .OE(N__2217),
            .DIN(N__2216),
            .DOUT(N__2215),
            .PACKAGEPIN(PMOD[22]));
    defparam PMOD_obuft_22_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_22_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_22_preio (
            .PADOEN(N__2217),
            .PADOUT(N__2216),
            .PADIN(N__2215),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_23_iopad (
            .OE(N__2208),
            .DIN(N__2207),
            .DOUT(N__2206),
            .PACKAGEPIN(PMOD[23]));
    defparam PMOD_obuft_23_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_23_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_23_preio (
            .PADOEN(N__2208),
            .PADOUT(N__2207),
            .PADIN(N__2206),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_24_iopad (
            .OE(N__2199),
            .DIN(N__2198),
            .DOUT(N__2197),
            .PACKAGEPIN(PMOD[24]));
    defparam PMOD_obuft_24_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_24_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_24_preio (
            .PADOEN(N__2199),
            .PADOUT(N__2198),
            .PADIN(N__2197),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_25_iopad (
            .OE(N__2190),
            .DIN(N__2189),
            .DOUT(N__2188),
            .PACKAGEPIN(PMOD[25]));
    defparam PMOD_obuft_25_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_25_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_25_preio (
            .PADOEN(N__2190),
            .PADOUT(N__2189),
            .PADIN(N__2188),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_26_iopad (
            .OE(N__2181),
            .DIN(N__2180),
            .DOUT(N__2179),
            .PACKAGEPIN(PMOD[26]));
    defparam PMOD_obuft_26_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_26_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_26_preio (
            .PADOEN(N__2181),
            .PADOUT(N__2180),
            .PADIN(N__2179),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_27_iopad (
            .OE(N__2172),
            .DIN(N__2171),
            .DOUT(N__2170),
            .PACKAGEPIN(PMOD[27]));
    defparam PMOD_obuft_27_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_27_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_27_preio (
            .PADOEN(N__2172),
            .PADOUT(N__2171),
            .PADIN(N__2170),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_28_iopad (
            .OE(N__2163),
            .DIN(N__2162),
            .DOUT(N__2161),
            .PACKAGEPIN(PMOD[28]));
    defparam PMOD_obuft_28_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_28_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_28_preio (
            .PADOEN(N__2163),
            .PADOUT(N__2162),
            .PADIN(N__2161),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_29_iopad (
            .OE(N__2154),
            .DIN(N__2153),
            .DOUT(N__2152),
            .PACKAGEPIN(PMOD[29]));
    defparam PMOD_obuft_29_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_29_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_29_preio (
            .PADOEN(N__2154),
            .PADOUT(N__2153),
            .PADIN(N__2152),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_3_iopad (
            .OE(N__2145),
            .DIN(N__2144),
            .DOUT(N__2143),
            .PACKAGEPIN(PMOD[3]));
    defparam PMOD_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_3_preio (
            .PADOEN(N__2145),
            .PADOUT(N__2144),
            .PADIN(N__2143),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_30_iopad (
            .OE(N__2136),
            .DIN(N__2135),
            .DOUT(N__2134),
            .PACKAGEPIN(PMOD[30]));
    defparam PMOD_obuft_30_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_30_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_30_preio (
            .PADOEN(N__2136),
            .PADOUT(N__2135),
            .PADIN(N__2134),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_31_iopad (
            .OE(N__2127),
            .DIN(N__2126),
            .DOUT(N__2125),
            .PACKAGEPIN(PMOD[31]));
    defparam PMOD_obuft_31_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_31_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_31_preio (
            .PADOEN(N__2127),
            .PADOUT(N__2126),
            .PADIN(N__2125),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_32_iopad (
            .OE(N__2118),
            .DIN(N__2117),
            .DOUT(N__2116),
            .PACKAGEPIN(PMOD[32]));
    defparam PMOD_obuft_32_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_32_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_32_preio (
            .PADOEN(N__2118),
            .PADOUT(N__2117),
            .PADIN(N__2116),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_33_iopad (
            .OE(N__2109),
            .DIN(N__2108),
            .DOUT(N__2107),
            .PACKAGEPIN(PMOD[33]));
    defparam PMOD_obuft_33_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_33_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_33_preio (
            .PADOEN(N__2109),
            .PADOUT(N__2108),
            .PADIN(N__2107),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_34_iopad (
            .OE(N__2100),
            .DIN(N__2099),
            .DOUT(N__2098),
            .PACKAGEPIN(PMOD[34]));
    defparam PMOD_obuft_34_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_34_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_34_preio (
            .PADOEN(N__2100),
            .PADOUT(N__2099),
            .PADIN(N__2098),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_35_iopad (
            .OE(N__2091),
            .DIN(N__2090),
            .DOUT(N__2089),
            .PACKAGEPIN(PMOD[35]));
    defparam PMOD_obuft_35_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_35_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_35_preio (
            .PADOEN(N__2091),
            .PADOUT(N__2090),
            .PADIN(N__2089),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_36_iopad (
            .OE(N__2082),
            .DIN(N__2081),
            .DOUT(N__2080),
            .PACKAGEPIN(PMOD[36]));
    defparam PMOD_obuft_36_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_36_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_36_preio (
            .PADOEN(N__2082),
            .PADOUT(N__2081),
            .PADIN(N__2080),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_37_iopad (
            .OE(N__2073),
            .DIN(N__2072),
            .DOUT(N__2071),
            .PACKAGEPIN(PMOD[37]));
    defparam PMOD_obuft_37_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_37_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_37_preio (
            .PADOEN(N__2073),
            .PADOUT(N__2072),
            .PADIN(N__2071),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_38_iopad (
            .OE(N__2064),
            .DIN(N__2063),
            .DOUT(N__2062),
            .PACKAGEPIN(PMOD[38]));
    defparam PMOD_obuft_38_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_38_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_38_preio (
            .PADOEN(N__2064),
            .PADOUT(N__2063),
            .PADIN(N__2062),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_39_iopad (
            .OE(N__2055),
            .DIN(N__2054),
            .DOUT(N__2053),
            .PACKAGEPIN(PMOD[39]));
    defparam PMOD_obuft_39_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_39_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_39_preio (
            .PADOEN(N__2055),
            .PADOUT(N__2054),
            .PADIN(N__2053),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_4_iopad (
            .OE(N__2046),
            .DIN(N__2045),
            .DOUT(N__2044),
            .PACKAGEPIN(PMOD[4]));
    defparam PMOD_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_4_preio (
            .PADOEN(N__2046),
            .PADOUT(N__2045),
            .PADIN(N__2044),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_40_iopad (
            .OE(N__2037),
            .DIN(N__2036),
            .DOUT(N__2035),
            .PACKAGEPIN(PMOD[40]));
    defparam PMOD_obuft_40_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_40_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_40_preio (
            .PADOEN(N__2037),
            .PADOUT(N__2036),
            .PADIN(N__2035),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_41_iopad (
            .OE(N__2028),
            .DIN(N__2027),
            .DOUT(N__2026),
            .PACKAGEPIN(PMOD[41]));
    defparam PMOD_obuft_41_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_41_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_41_preio (
            .PADOEN(N__2028),
            .PADOUT(N__2027),
            .PADIN(N__2026),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_42_iopad (
            .OE(N__2019),
            .DIN(N__2018),
            .DOUT(N__2017),
            .PACKAGEPIN(PMOD[42]));
    defparam PMOD_obuft_42_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_42_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_42_preio (
            .PADOEN(N__2019),
            .PADOUT(N__2018),
            .PADIN(N__2017),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_43_iopad (
            .OE(N__2010),
            .DIN(N__2009),
            .DOUT(N__2008),
            .PACKAGEPIN(PMOD[43]));
    defparam PMOD_obuft_43_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_43_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_43_preio (
            .PADOEN(N__2010),
            .PADOUT(N__2009),
            .PADIN(N__2008),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_44_iopad (
            .OE(N__2001),
            .DIN(N__2000),
            .DOUT(N__1999),
            .PACKAGEPIN(PMOD[44]));
    defparam PMOD_obuft_44_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_44_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_44_preio (
            .PADOEN(N__2001),
            .PADOUT(N__2000),
            .PADIN(N__1999),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_45_iopad (
            .OE(N__1992),
            .DIN(N__1991),
            .DOUT(N__1990),
            .PACKAGEPIN(PMOD[45]));
    defparam PMOD_obuft_45_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_45_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_45_preio (
            .PADOEN(N__1992),
            .PADOUT(N__1991),
            .PADIN(N__1990),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_46_iopad (
            .OE(N__1983),
            .DIN(N__1982),
            .DOUT(N__1981),
            .PACKAGEPIN(PMOD[46]));
    defparam PMOD_obuft_46_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_46_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_46_preio (
            .PADOEN(N__1983),
            .PADOUT(N__1982),
            .PADIN(N__1981),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_47_iopad (
            .OE(N__1974),
            .DIN(N__1973),
            .DOUT(N__1972),
            .PACKAGEPIN(PMOD[47]));
    defparam PMOD_obuft_47_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_47_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_47_preio (
            .PADOEN(N__1974),
            .PADOUT(N__1973),
            .PADIN(N__1972),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_48_iopad (
            .OE(N__1965),
            .DIN(N__1964),
            .DOUT(N__1963),
            .PACKAGEPIN(PMOD[48]));
    defparam PMOD_obuft_48_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_48_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_48_preio (
            .PADOEN(N__1965),
            .PADOUT(N__1964),
            .PADIN(N__1963),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_49_iopad (
            .OE(N__1956),
            .DIN(N__1955),
            .DOUT(N__1954),
            .PACKAGEPIN(PMOD[49]));
    defparam PMOD_obuft_49_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_49_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_49_preio (
            .PADOEN(N__1956),
            .PADOUT(N__1955),
            .PADIN(N__1954),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_5_iopad (
            .OE(N__1947),
            .DIN(N__1946),
            .DOUT(N__1945),
            .PACKAGEPIN(PMOD[5]));
    defparam PMOD_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_5_preio (
            .PADOEN(N__1947),
            .PADOUT(N__1946),
            .PADIN(N__1945),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_50_iopad (
            .OE(N__1938),
            .DIN(N__1937),
            .DOUT(N__1936),
            .PACKAGEPIN(PMOD[50]));
    defparam PMOD_obuft_50_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_50_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_50_preio (
            .PADOEN(N__1938),
            .PADOUT(N__1937),
            .PADIN(N__1936),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_51_iopad (
            .OE(N__1929),
            .DIN(N__1928),
            .DOUT(N__1927),
            .PACKAGEPIN(PMOD[51]));
    defparam PMOD_obuft_51_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_51_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_51_preio (
            .PADOEN(N__1929),
            .PADOUT(N__1928),
            .PADIN(N__1927),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_6_iopad (
            .OE(N__1920),
            .DIN(N__1919),
            .DOUT(N__1918),
            .PACKAGEPIN(PMOD[6]));
    defparam PMOD_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_6_preio (
            .PADOEN(N__1920),
            .PADOUT(N__1919),
            .PADIN(N__1918),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_7_iopad (
            .OE(N__1911),
            .DIN(N__1910),
            .DOUT(N__1909),
            .PACKAGEPIN(PMOD[7]));
    defparam PMOD_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_7_preio (
            .PADOEN(N__1911),
            .PADOUT(N__1910),
            .PADIN(N__1909),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_8_iopad (
            .OE(N__1902),
            .DIN(N__1901),
            .DOUT(N__1900),
            .PACKAGEPIN(PMOD[8]));
    defparam PMOD_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_8_preio (
            .PADOEN(N__1902),
            .PADOUT(N__1901),
            .PADIN(N__1900),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PMOD_obuft_9_iopad (
            .OE(N__1893),
            .DIN(N__1892),
            .DOUT(N__1891),
            .PACKAGEPIN(PMOD[9]));
    defparam PMOD_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam PMOD_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO PMOD_obuft_9_preio (
            .PADOEN(N__1893),
            .PADOUT(N__1892),
            .PADIN(N__1891),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD RAMCS_obuf_iopad (
            .OE(N__1884),
            .DIN(N__1883),
            .DOUT(N__1882),
            .PACKAGEPIN(RAMCS));
    defparam RAMCS_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMCS_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMCS_obuf_preio (
            .PADOEN(N__1884),
            .PADOUT(N__1883),
            .PADIN(N__1882),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1469),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD RAMOE_obuf_iopad (
            .OE(N__1875),
            .DIN(N__1874),
            .DOUT(N__1873),
            .PACKAGEPIN(RAMOE));
    defparam RAMOE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMOE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMOE_obuf_preio (
            .PADOEN(N__1875),
            .PADOUT(N__1874),
            .PADIN(N__1873),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1458),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD RAMWE_obuf_iopad (
            .OE(N__1866),
            .DIN(N__1865),
            .DOUT(N__1864),
            .PACKAGEPIN(RAMWE));
    defparam RAMWE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMWE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMWE_obuf_preio (
            .PADOEN(N__1866),
            .PADOUT(N__1865),
            .PADIN(N__1864),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1468),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__273 (
            .O(N__1847),
            .I(N__1843));
    IoInMux I__272 (
            .O(N__1846),
            .I(N__1840));
    LocalMux I__271 (
            .O(N__1843),
            .I(N__1835));
    LocalMux I__270 (
            .O(N__1840),
            .I(N__1835));
    IoSpan4Mux I__269 (
            .O(N__1835),
            .I(N__1832));
    Span4Mux_s2_v I__268 (
            .O(N__1832),
            .I(N__1828));
    InMux I__267 (
            .O(N__1831),
            .I(N__1825));
    Span4Mux_v I__266 (
            .O(N__1828),
            .I(N__1820));
    LocalMux I__265 (
            .O(N__1825),
            .I(N__1820));
    Span4Mux_h I__264 (
            .O(N__1820),
            .I(N__1817));
    Span4Mux_v I__263 (
            .O(N__1817),
            .I(N__1813));
    InMux I__262 (
            .O(N__1816),
            .I(N__1810));
    Odrv4 I__261 (
            .O(N__1813),
            .I(PMOD_c_52));
    LocalMux I__260 (
            .O(N__1810),
            .I(PMOD_c_52));
    IoInMux I__259 (
            .O(N__1805),
            .I(N__1802));
    LocalMux I__258 (
            .O(N__1802),
            .I(N__1798));
    IoInMux I__257 (
            .O(N__1801),
            .I(N__1795));
    IoSpan4Mux I__256 (
            .O(N__1798),
            .I(N__1792));
    LocalMux I__255 (
            .O(N__1795),
            .I(N__1789));
    Span4Mux_s2_h I__254 (
            .O(N__1792),
            .I(N__1784));
    Span4Mux_s2_v I__253 (
            .O(N__1789),
            .I(N__1784));
    Span4Mux_v I__252 (
            .O(N__1784),
            .I(N__1781));
    Odrv4 I__251 (
            .O(N__1781),
            .I(PMOD_c_i_52));
    CascadeMux I__250 (
            .O(N__1778),
            .I(N__1775));
    InMux I__249 (
            .O(N__1775),
            .I(N__1772));
    LocalMux I__248 (
            .O(N__1772),
            .I(\my_alternate.countZ0Z_17 ));
    InMux I__247 (
            .O(N__1769),
            .I(\my_alternate.count_cry_16 ));
    CascadeMux I__246 (
            .O(N__1766),
            .I(N__1763));
    InMux I__245 (
            .O(N__1763),
            .I(N__1760));
    LocalMux I__244 (
            .O(N__1760),
            .I(\my_alternate.countZ0Z_18 ));
    InMux I__243 (
            .O(N__1757),
            .I(\my_alternate.count_cry_17 ));
    CascadeMux I__242 (
            .O(N__1754),
            .I(N__1751));
    InMux I__241 (
            .O(N__1751),
            .I(N__1748));
    LocalMux I__240 (
            .O(N__1748),
            .I(\my_alternate.countZ0Z_19 ));
    InMux I__239 (
            .O(N__1745),
            .I(\my_alternate.count_cry_18 ));
    CascadeMux I__238 (
            .O(N__1742),
            .I(N__1739));
    InMux I__237 (
            .O(N__1739),
            .I(N__1736));
    LocalMux I__236 (
            .O(N__1736),
            .I(\my_alternate.countZ0Z_20 ));
    InMux I__235 (
            .O(N__1733),
            .I(\my_alternate.count_cry_19 ));
    CascadeMux I__234 (
            .O(N__1730),
            .I(N__1727));
    InMux I__233 (
            .O(N__1727),
            .I(N__1724));
    LocalMux I__232 (
            .O(N__1724),
            .I(\my_alternate.countZ0Z_21 ));
    InMux I__231 (
            .O(N__1721),
            .I(\my_alternate.count_cry_20 ));
    CascadeMux I__230 (
            .O(N__1718),
            .I(N__1715));
    InMux I__229 (
            .O(N__1715),
            .I(N__1712));
    LocalMux I__228 (
            .O(N__1712),
            .I(\my_alternate.countZ0Z_22 ));
    InMux I__227 (
            .O(N__1709),
            .I(\my_alternate.count_cry_21 ));
    CascadeMux I__226 (
            .O(N__1706),
            .I(N__1703));
    InMux I__225 (
            .O(N__1703),
            .I(N__1700));
    LocalMux I__224 (
            .O(N__1700),
            .I(\my_alternate.countZ0Z_23 ));
    InMux I__223 (
            .O(N__1697),
            .I(\my_alternate.count_cry_22 ));
    InMux I__222 (
            .O(N__1694),
            .I(bfn_19_9_0_));
    ClkMux I__221 (
            .O(N__1691),
            .I(N__1679));
    ClkMux I__220 (
            .O(N__1690),
            .I(N__1679));
    ClkMux I__219 (
            .O(N__1689),
            .I(N__1679));
    ClkMux I__218 (
            .O(N__1688),
            .I(N__1679));
    GlobalMux I__217 (
            .O(N__1679),
            .I(N__1676));
    gio2CtrlBuf I__216 (
            .O(N__1676),
            .I(clk_c_g));
    CascadeMux I__215 (
            .O(N__1673),
            .I(N__1670));
    InMux I__214 (
            .O(N__1670),
            .I(N__1667));
    LocalMux I__213 (
            .O(N__1667),
            .I(\my_alternate.countZ0Z_9 ));
    InMux I__212 (
            .O(N__1664),
            .I(\my_alternate.count_cry_8 ));
    CascadeMux I__211 (
            .O(N__1661),
            .I(N__1658));
    InMux I__210 (
            .O(N__1658),
            .I(N__1655));
    LocalMux I__209 (
            .O(N__1655),
            .I(\my_alternate.countZ0Z_10 ));
    InMux I__208 (
            .O(N__1652),
            .I(\my_alternate.count_cry_9 ));
    CascadeMux I__207 (
            .O(N__1649),
            .I(N__1646));
    InMux I__206 (
            .O(N__1646),
            .I(N__1643));
    LocalMux I__205 (
            .O(N__1643),
            .I(\my_alternate.countZ0Z_11 ));
    InMux I__204 (
            .O(N__1640),
            .I(\my_alternate.count_cry_10 ));
    CascadeMux I__203 (
            .O(N__1637),
            .I(N__1634));
    InMux I__202 (
            .O(N__1634),
            .I(N__1631));
    LocalMux I__201 (
            .O(N__1631),
            .I(\my_alternate.countZ0Z_12 ));
    InMux I__200 (
            .O(N__1628),
            .I(\my_alternate.count_cry_11 ));
    CascadeMux I__199 (
            .O(N__1625),
            .I(N__1622));
    InMux I__198 (
            .O(N__1622),
            .I(N__1619));
    LocalMux I__197 (
            .O(N__1619),
            .I(\my_alternate.countZ0Z_13 ));
    InMux I__196 (
            .O(N__1616),
            .I(\my_alternate.count_cry_12 ));
    CascadeMux I__195 (
            .O(N__1613),
            .I(N__1610));
    InMux I__194 (
            .O(N__1610),
            .I(N__1607));
    LocalMux I__193 (
            .O(N__1607),
            .I(\my_alternate.countZ0Z_14 ));
    InMux I__192 (
            .O(N__1604),
            .I(\my_alternate.count_cry_13 ));
    CascadeMux I__191 (
            .O(N__1601),
            .I(N__1598));
    InMux I__190 (
            .O(N__1598),
            .I(N__1595));
    LocalMux I__189 (
            .O(N__1595),
            .I(\my_alternate.countZ0Z_15 ));
    InMux I__188 (
            .O(N__1592),
            .I(\my_alternate.count_cry_14 ));
    CascadeMux I__187 (
            .O(N__1589),
            .I(N__1586));
    InMux I__186 (
            .O(N__1586),
            .I(N__1583));
    LocalMux I__185 (
            .O(N__1583),
            .I(\my_alternate.countZ0Z_16 ));
    InMux I__184 (
            .O(N__1580),
            .I(bfn_19_8_0_));
    CascadeMux I__183 (
            .O(N__1577),
            .I(N__1574));
    InMux I__182 (
            .O(N__1574),
            .I(N__1571));
    LocalMux I__181 (
            .O(N__1571),
            .I(\my_alternate.countZ0Z_0 ));
    InMux I__180 (
            .O(N__1568),
            .I(bfn_19_6_0_));
    CascadeMux I__179 (
            .O(N__1565),
            .I(N__1562));
    InMux I__178 (
            .O(N__1562),
            .I(N__1559));
    LocalMux I__177 (
            .O(N__1559),
            .I(\my_alternate.countZ0Z_1 ));
    InMux I__176 (
            .O(N__1556),
            .I(\my_alternate.count_cry_0 ));
    CascadeMux I__175 (
            .O(N__1553),
            .I(N__1550));
    InMux I__174 (
            .O(N__1550),
            .I(N__1547));
    LocalMux I__173 (
            .O(N__1547),
            .I(\my_alternate.countZ0Z_2 ));
    InMux I__172 (
            .O(N__1544),
            .I(\my_alternate.count_cry_1 ));
    CascadeMux I__171 (
            .O(N__1541),
            .I(N__1538));
    InMux I__170 (
            .O(N__1538),
            .I(N__1535));
    LocalMux I__169 (
            .O(N__1535),
            .I(\my_alternate.countZ0Z_3 ));
    InMux I__168 (
            .O(N__1532),
            .I(\my_alternate.count_cry_2 ));
    CascadeMux I__167 (
            .O(N__1529),
            .I(N__1526));
    InMux I__166 (
            .O(N__1526),
            .I(N__1523));
    LocalMux I__165 (
            .O(N__1523),
            .I(\my_alternate.countZ0Z_4 ));
    InMux I__164 (
            .O(N__1520),
            .I(\my_alternate.count_cry_3 ));
    CascadeMux I__163 (
            .O(N__1517),
            .I(N__1514));
    InMux I__162 (
            .O(N__1514),
            .I(N__1511));
    LocalMux I__161 (
            .O(N__1511),
            .I(\my_alternate.countZ0Z_5 ));
    InMux I__160 (
            .O(N__1508),
            .I(\my_alternate.count_cry_4 ));
    CascadeMux I__159 (
            .O(N__1505),
            .I(N__1502));
    InMux I__158 (
            .O(N__1502),
            .I(N__1499));
    LocalMux I__157 (
            .O(N__1499),
            .I(\my_alternate.countZ0Z_6 ));
    InMux I__156 (
            .O(N__1496),
            .I(\my_alternate.count_cry_5 ));
    CascadeMux I__155 (
            .O(N__1493),
            .I(N__1490));
    InMux I__154 (
            .O(N__1490),
            .I(N__1487));
    LocalMux I__153 (
            .O(N__1487),
            .I(\my_alternate.countZ0Z_7 ));
    InMux I__152 (
            .O(N__1484),
            .I(\my_alternate.count_cry_6 ));
    CascadeMux I__151 (
            .O(N__1481),
            .I(N__1478));
    InMux I__150 (
            .O(N__1478),
            .I(N__1475));
    LocalMux I__149 (
            .O(N__1475),
            .I(\my_alternate.countZ0Z_8 ));
    InMux I__148 (
            .O(N__1472),
            .I(bfn_19_7_0_));
    IoInMux I__147 (
            .O(N__1469),
            .I(N__1465));
    IoInMux I__146 (
            .O(N__1468),
            .I(N__1462));
    LocalMux I__145 (
            .O(N__1465),
            .I(N__1459));
    LocalMux I__144 (
            .O(N__1462),
            .I(N__1455));
    Span4Mux_s2_v I__143 (
            .O(N__1459),
            .I(N__1452));
    IoInMux I__142 (
            .O(N__1458),
            .I(N__1449));
    Span4Mux_s3_v I__141 (
            .O(N__1455),
            .I(N__1446));
    Sp12to4 I__140 (
            .O(N__1452),
            .I(N__1443));
    LocalMux I__139 (
            .O(N__1449),
            .I(N__1440));
    Span4Mux_h I__138 (
            .O(N__1446),
            .I(N__1437));
    Span12Mux_h I__137 (
            .O(N__1443),
            .I(N__1434));
    Span12Mux_s5_v I__136 (
            .O(N__1440),
            .I(N__1431));
    Span4Mux_v I__135 (
            .O(N__1437),
            .I(N__1428));
    Span12Mux_v I__134 (
            .O(N__1434),
            .I(N__1425));
    Span12Mux_v I__133 (
            .O(N__1431),
            .I(N__1422));
    Span4Mux_v I__132 (
            .O(N__1428),
            .I(N__1419));
    Odrv12 I__131 (
            .O(N__1425),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__130 (
            .O(N__1422),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__129 (
            .O(N__1419),
            .I(CONSTANT_ONE_NET));
    defparam IN_MUX_bfv_19_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_6_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(\my_alternate.count_cry_7 ),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_19_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_8_0_ (
            .carryinitin(\my_alternate.count_cry_15 ),
            .carryinitout(bfn_19_8_0_));
    defparam IN_MUX_bfv_19_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_9_0_ (
            .carryinitin(\my_alternate.count_cry_23 ),
            .carryinitout(bfn_19_9_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_18_12_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_18_12_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_18_12_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_18_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_0_LC_19_6_0 .C_ON=1'b1;
    defparam \my_alternate.count_0_LC_19_6_0 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_0_LC_19_6_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_0_LC_19_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1577),
            .in3(N__1568),
            .lcout(\my_alternate.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_19_6_0_),
            .carryout(\my_alternate.count_cry_0 ),
            .clk(N__1691),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_1_LC_19_6_1 .C_ON=1'b1;
    defparam \my_alternate.count_1_LC_19_6_1 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_1_LC_19_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_1_LC_19_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1565),
            .in3(N__1556),
            .lcout(\my_alternate.countZ0Z_1 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_0 ),
            .carryout(\my_alternate.count_cry_1 ),
            .clk(N__1691),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_2_LC_19_6_2 .C_ON=1'b1;
    defparam \my_alternate.count_2_LC_19_6_2 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_2_LC_19_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_2_LC_19_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1553),
            .in3(N__1544),
            .lcout(\my_alternate.countZ0Z_2 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_1 ),
            .carryout(\my_alternate.count_cry_2 ),
            .clk(N__1691),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_3_LC_19_6_3 .C_ON=1'b1;
    defparam \my_alternate.count_3_LC_19_6_3 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_3_LC_19_6_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_3_LC_19_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1541),
            .in3(N__1532),
            .lcout(\my_alternate.countZ0Z_3 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_2 ),
            .carryout(\my_alternate.count_cry_3 ),
            .clk(N__1691),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_4_LC_19_6_4 .C_ON=1'b1;
    defparam \my_alternate.count_4_LC_19_6_4 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_4_LC_19_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_4_LC_19_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1529),
            .in3(N__1520),
            .lcout(\my_alternate.countZ0Z_4 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_3 ),
            .carryout(\my_alternate.count_cry_4 ),
            .clk(N__1691),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_5_LC_19_6_5 .C_ON=1'b1;
    defparam \my_alternate.count_5_LC_19_6_5 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_5_LC_19_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_5_LC_19_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1517),
            .in3(N__1508),
            .lcout(\my_alternate.countZ0Z_5 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_4 ),
            .carryout(\my_alternate.count_cry_5 ),
            .clk(N__1691),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_6_LC_19_6_6 .C_ON=1'b1;
    defparam \my_alternate.count_6_LC_19_6_6 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_6_LC_19_6_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_6_LC_19_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1505),
            .in3(N__1496),
            .lcout(\my_alternate.countZ0Z_6 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_5 ),
            .carryout(\my_alternate.count_cry_6 ),
            .clk(N__1691),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_7_LC_19_6_7 .C_ON=1'b1;
    defparam \my_alternate.count_7_LC_19_6_7 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_7_LC_19_6_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_7_LC_19_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1493),
            .in3(N__1484),
            .lcout(\my_alternate.countZ0Z_7 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_6 ),
            .carryout(\my_alternate.count_cry_7 ),
            .clk(N__1691),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_8_LC_19_7_0 .C_ON=1'b1;
    defparam \my_alternate.count_8_LC_19_7_0 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_8_LC_19_7_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_8_LC_19_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1481),
            .in3(N__1472),
            .lcout(\my_alternate.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(\my_alternate.count_cry_8 ),
            .clk(N__1690),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_9_LC_19_7_1 .C_ON=1'b1;
    defparam \my_alternate.count_9_LC_19_7_1 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_9_LC_19_7_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_9_LC_19_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1673),
            .in3(N__1664),
            .lcout(\my_alternate.countZ0Z_9 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_8 ),
            .carryout(\my_alternate.count_cry_9 ),
            .clk(N__1690),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_10_LC_19_7_2 .C_ON=1'b1;
    defparam \my_alternate.count_10_LC_19_7_2 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_10_LC_19_7_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_10_LC_19_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1661),
            .in3(N__1652),
            .lcout(\my_alternate.countZ0Z_10 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_9 ),
            .carryout(\my_alternate.count_cry_10 ),
            .clk(N__1690),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_11_LC_19_7_3 .C_ON=1'b1;
    defparam \my_alternate.count_11_LC_19_7_3 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_11_LC_19_7_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_11_LC_19_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1649),
            .in3(N__1640),
            .lcout(\my_alternate.countZ0Z_11 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_10 ),
            .carryout(\my_alternate.count_cry_11 ),
            .clk(N__1690),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_12_LC_19_7_4 .C_ON=1'b1;
    defparam \my_alternate.count_12_LC_19_7_4 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_12_LC_19_7_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_12_LC_19_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1637),
            .in3(N__1628),
            .lcout(\my_alternate.countZ0Z_12 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_11 ),
            .carryout(\my_alternate.count_cry_12 ),
            .clk(N__1690),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_13_LC_19_7_5 .C_ON=1'b1;
    defparam \my_alternate.count_13_LC_19_7_5 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_13_LC_19_7_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_13_LC_19_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1625),
            .in3(N__1616),
            .lcout(\my_alternate.countZ0Z_13 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_12 ),
            .carryout(\my_alternate.count_cry_13 ),
            .clk(N__1690),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_14_LC_19_7_6 .C_ON=1'b1;
    defparam \my_alternate.count_14_LC_19_7_6 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_14_LC_19_7_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_14_LC_19_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1613),
            .in3(N__1604),
            .lcout(\my_alternate.countZ0Z_14 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_13 ),
            .carryout(\my_alternate.count_cry_14 ),
            .clk(N__1690),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_15_LC_19_7_7 .C_ON=1'b1;
    defparam \my_alternate.count_15_LC_19_7_7 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_15_LC_19_7_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_15_LC_19_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1601),
            .in3(N__1592),
            .lcout(\my_alternate.countZ0Z_15 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_14 ),
            .carryout(\my_alternate.count_cry_15 ),
            .clk(N__1690),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_16_LC_19_8_0 .C_ON=1'b1;
    defparam \my_alternate.count_16_LC_19_8_0 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_16_LC_19_8_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_16_LC_19_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1589),
            .in3(N__1580),
            .lcout(\my_alternate.countZ0Z_16 ),
            .ltout(),
            .carryin(bfn_19_8_0_),
            .carryout(\my_alternate.count_cry_16 ),
            .clk(N__1689),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_17_LC_19_8_1 .C_ON=1'b1;
    defparam \my_alternate.count_17_LC_19_8_1 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_17_LC_19_8_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_17_LC_19_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1778),
            .in3(N__1769),
            .lcout(\my_alternate.countZ0Z_17 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_16 ),
            .carryout(\my_alternate.count_cry_17 ),
            .clk(N__1689),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_18_LC_19_8_2 .C_ON=1'b1;
    defparam \my_alternate.count_18_LC_19_8_2 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_18_LC_19_8_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_18_LC_19_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1766),
            .in3(N__1757),
            .lcout(\my_alternate.countZ0Z_18 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_17 ),
            .carryout(\my_alternate.count_cry_18 ),
            .clk(N__1689),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_19_LC_19_8_3 .C_ON=1'b1;
    defparam \my_alternate.count_19_LC_19_8_3 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_19_LC_19_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_19_LC_19_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1754),
            .in3(N__1745),
            .lcout(\my_alternate.countZ0Z_19 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_18 ),
            .carryout(\my_alternate.count_cry_19 ),
            .clk(N__1689),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_20_LC_19_8_4 .C_ON=1'b1;
    defparam \my_alternate.count_20_LC_19_8_4 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_20_LC_19_8_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_20_LC_19_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1742),
            .in3(N__1733),
            .lcout(\my_alternate.countZ0Z_20 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_19 ),
            .carryout(\my_alternate.count_cry_20 ),
            .clk(N__1689),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_21_LC_19_8_5 .C_ON=1'b1;
    defparam \my_alternate.count_21_LC_19_8_5 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_21_LC_19_8_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_21_LC_19_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1730),
            .in3(N__1721),
            .lcout(\my_alternate.countZ0Z_21 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_20 ),
            .carryout(\my_alternate.count_cry_21 ),
            .clk(N__1689),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_22_LC_19_8_6 .C_ON=1'b1;
    defparam \my_alternate.count_22_LC_19_8_6 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_22_LC_19_8_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_22_LC_19_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1718),
            .in3(N__1709),
            .lcout(\my_alternate.countZ0Z_22 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_21 ),
            .carryout(\my_alternate.count_cry_22 ),
            .clk(N__1689),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_23_LC_19_8_7 .C_ON=1'b1;
    defparam \my_alternate.count_23_LC_19_8_7 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_23_LC_19_8_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \my_alternate.count_23_LC_19_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1706),
            .in3(N__1697),
            .lcout(\my_alternate.countZ0Z_23 ),
            .ltout(),
            .carryin(\my_alternate.count_cry_22 ),
            .carryout(\my_alternate.count_cry_23 ),
            .clk(N__1689),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_24_LC_19_9_0 .C_ON=1'b0;
    defparam \my_alternate.count_24_LC_19_9_0 .SEQ_MODE=4'b1000;
    defparam \my_alternate.count_24_LC_19_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \my_alternate.count_24_LC_19_9_0  (
            .in0(_gnd_net_),
            .in1(N__1816),
            .in2(_gnd_net_),
            .in3(N__1694),
            .lcout(PMOD_c_52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1688),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_alternate.count_RNIQ674_24_LC_23_1_1 .C_ON=1'b0;
    defparam \my_alternate.count_RNIQ674_24_LC_23_1_1 .SEQ_MODE=4'b0000;
    defparam \my_alternate.count_RNIQ674_24_LC_23_1_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \my_alternate.count_RNIQ674_24_LC_23_1_1  (
            .in0(N__1831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PMOD_c_i_52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // chip
